module CPU(
    input logic clk,
    input logic n_reset,
    input logic [3:0] addr,
    input logic [7:0] data,
    input logic [3:0] switch,
    input logic [3:0] switch,
)
